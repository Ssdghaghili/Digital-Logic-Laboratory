module mux8(sel,in1,in2,out);
  input sel;
  input [7:0] in1;
  input [7:0] in2;
  output [7:0] out;
  assign out = sel?in1:in2;
endmodule
      
  
