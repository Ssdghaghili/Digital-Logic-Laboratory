module shr2bit(serIn , shen , clk,rst,clkEn,portnum);
  input serIn,shen,clk,rst,clkEn;
  output[1:0] portnum;
  reg [1:0] shift;
  always@(posedge clkEn , posedge rst)
  begin
    if(rst)
      shift <= 2'b0;
    else if(shen)
      shift <= {shift[0] , serIn};
  end
  assign portnum=shift;
endmodule
